module data_cache #(
    parameter XLEN = 32
) (
    input  logic clk,
    input  logic rst,
    input  logic [XLEN-1:0] A,
    input  logic [XLEN-1:0] WD,
    input  logic WE,
    input  logic [31:0] mem_rd_data, // data read from main mem
    output logic [31:0] cache_dout // data out to cpu
);

logic [20:0] tag;
logic [8:0] set;

// WAY 0 ARRAYS
logic        v_way0    [511:0]; // valid bit
logic        d_way0    [511:0]; // dirty bit
logic [20:0] tag_way0  [511:0]; // tag
logic [31:0] data_way0 [511:0]; // data
// WAY 1 ARRAYS
logic        v_way1    [511:0]; // valid bit
logic        d_way1    [511:0]; // dirty bit
logic [20:0] tag_way1  [511:0]; // tag
logic [31:0] data_way1 [511:0]; // data

logic u_bit [511:0]; // 0 = way0 accessed most recently, 1 = way1 accessed most recently

logic hit0; // way 0 hit
logic hit1; // way 1 hit
logic hit;

logic [31:0] mem_rd_data;
//logic [31:0] ram_write;
//logic ram_write_en;

// clear cache valid bits on startup
initial begin
    for (int i = 0; i < 512; i++) begin
        v_way0[i] = 0;
        v_way1[i] = 0;
        u_bit [i] = 0;
        d_way0[i] = 0;
        d_way1[i] = 0;
    end
end

assign tag = A[31:11];
assign set = A[10:2];

assign hit0 = v_way0[set] && (tag_way0[set] == tag);
assign hit1 = v_way1[set] && (tag_way1[set] == tag);
assign hit  = hit0 || hit1;

always_comb begin
    if (hit0)      cache_dout = data_way0[set];
    else if (hit1) cache_dout = data_way1[set];
    else           cache_dout = mem_rd_data;
end

always_ff @(posedge clk) begin
    // reset valid bits on a rst signal
    if (rst) begin
        for(int i=0; i<512; i++) begin
            v_way0[i] = 0;
            v_way1[i] = 0;
            u_bit [i] = 0;
            d_way0[i] = 0;
            d_way1[i] = 0;
        end
    end
    else begin
        // write: on a hit write to cache and set dirty bit true 
        if (WE) begin
            if (hit0) begin
                data_way0[set] <= WD;
                u_bit[set]  <= 0;
                d_way0[set] <= 1;
            end
            else if (hit1) begin
                data_way1[set] <= WD;
                u_bit[set]  <= 1;
                d_way1[set] <= 1;
            end
        end
        // on a read miss, bring data from ram to cache
        else if (!hit && !WE) begin
            ram_write_en <= 0;
            if (u_bit[set] == 1) begin // 1 most recently used so load into 0

                // if(d_way0[set] == 1) begin // write data from cache to memory before getting evicted 
                //     ram_write_en <= 1;
                //     ram_write <= data_way0[set];
                // end
                
                data_way0[set] <= mem_rd_data;
                tag_way0[set]  <= tag;
                v_way0[set] <= 1;
                d_way0[set] <= 0;
                u_bit[set]  <= 0; // way 0 most recently used
            end
            else begin // 0 most recently used so load into 1

                // if(d_way1[set] == 1) begin // write data from cache to memory before getting evicted 
                //     ram_write_en <= 1;
                //     ram_write <= data_way1[set];
                // end

                data_way1[set] <= mem_rd_data;
                tag_way1[set]  <= tag;
                v_way1[set] <= 1;
                d_way1[set] <= 0;
                u_bit[set]  <= 1; // way 1 most recently used
            end
        end
        else if (hit && !WE) begin // read hit: update
            if (hit0) u_bit[set] <= 1;
            if (hit1) u_bit[set] <= 0;
        end
    end
end

endmodule
